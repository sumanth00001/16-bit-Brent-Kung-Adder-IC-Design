magic
tech sky130A
magscale 1 2
timestamp 1668419820
<< nwell >>
rect 1066 116677 178886 117243
rect 1066 115589 178886 116155
rect 1066 114501 178886 115067
rect 1066 113413 178886 113979
rect 1066 112325 178886 112891
rect 1066 111237 178886 111803
rect 1066 110149 178886 110715
rect 1066 109061 178886 109627
rect 1066 107973 178886 108539
rect 1066 106885 178886 107451
rect 1066 105797 178886 106363
rect 1066 104709 178886 105275
rect 1066 103621 178886 104187
rect 1066 102533 178886 103099
rect 1066 101445 178886 102011
rect 1066 100357 178886 100923
rect 1066 99269 178886 99835
rect 1066 98181 178886 98747
rect 1066 97093 178886 97659
rect 1066 96005 178886 96571
rect 1066 94917 178886 95483
rect 1066 93829 178886 94395
rect 1066 92741 178886 93307
rect 1066 91653 178886 92219
rect 1066 90565 178886 91131
rect 1066 89477 178886 90043
rect 1066 88389 178886 88955
rect 1066 87301 178886 87867
rect 1066 86213 178886 86779
rect 1066 85125 178886 85691
rect 1066 84037 178886 84603
rect 1066 82949 178886 83515
rect 1066 81861 178886 82427
rect 1066 80773 178886 81339
rect 1066 79685 178886 80251
rect 1066 78597 178886 79163
rect 1066 77509 178886 78075
rect 1066 76421 178886 76987
rect 1066 75333 178886 75899
rect 1066 74245 178886 74811
rect 1066 73157 178886 73723
rect 1066 72069 178886 72635
rect 1066 70981 178886 71547
rect 1066 69893 178886 70459
rect 1066 68805 178886 69371
rect 1066 67717 178886 68283
rect 1066 66629 178886 67195
rect 1066 65541 178886 66107
rect 1066 64453 178886 65019
rect 1066 63365 178886 63931
rect 1066 62277 178886 62843
rect 1066 61189 178886 61755
rect 1066 60101 178886 60667
rect 1066 59013 178886 59579
rect 1066 57925 178886 58491
rect 1066 56837 178886 57403
rect 1066 55749 178886 56315
rect 1066 54661 178886 55227
rect 1066 53573 178886 54139
rect 1066 52485 178886 53051
rect 1066 51397 178886 51963
rect 1066 50309 178886 50875
rect 1066 49221 178886 49787
rect 1066 48133 178886 48699
rect 1066 47045 178886 47611
rect 1066 45957 178886 46523
rect 1066 44869 178886 45435
rect 1066 43781 178886 44347
rect 1066 42693 178886 43259
rect 1066 41605 178886 42171
rect 1066 40517 178886 41083
rect 1066 39429 178886 39995
rect 1066 38341 178886 38907
rect 1066 37253 178886 37819
rect 1066 36165 178886 36731
rect 1066 35077 178886 35643
rect 1066 33989 178886 34555
rect 1066 32901 178886 33467
rect 1066 31813 178886 32379
rect 1066 30725 178886 31291
rect 1066 29637 178886 30203
rect 1066 28549 178886 29115
rect 1066 27461 178886 28027
rect 1066 26373 178886 26939
rect 1066 25285 178886 25851
rect 1066 24197 178886 24763
rect 1066 23109 178886 23675
rect 1066 22021 178886 22587
rect 1066 20933 178886 21499
rect 1066 19845 178886 20411
rect 1066 18757 178886 19323
rect 1066 17669 178886 18235
rect 1066 16581 178886 17147
rect 1066 15493 178886 16059
rect 1066 14405 178886 14971
rect 1066 13317 178886 13883
rect 1066 12229 178886 12795
rect 1066 11141 178886 11707
rect 1066 10053 178886 10619
rect 1066 8965 178886 9531
rect 1066 7877 178886 8443
rect 1066 6789 178886 7355
rect 1066 5701 178886 6267
rect 1066 4613 178886 5179
rect 1066 3525 178886 4091
rect 1066 2437 178886 3003
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 2128 178848 117552
<< metal2 >>
rect 1582 119200 1638 120000
rect 3146 119200 3202 120000
rect 4710 119200 4766 120000
rect 6274 119200 6330 120000
rect 7838 119200 7894 120000
rect 9402 119200 9458 120000
rect 10966 119200 11022 120000
rect 12530 119200 12586 120000
rect 14094 119200 14150 120000
rect 15658 119200 15714 120000
rect 17222 119200 17278 120000
rect 18786 119200 18842 120000
rect 20350 119200 20406 120000
rect 21914 119200 21970 120000
rect 23478 119200 23534 120000
rect 25042 119200 25098 120000
rect 26606 119200 26662 120000
rect 28170 119200 28226 120000
rect 29734 119200 29790 120000
rect 31298 119200 31354 120000
rect 32862 119200 32918 120000
rect 34426 119200 34482 120000
rect 35990 119200 36046 120000
rect 37554 119200 37610 120000
rect 39118 119200 39174 120000
rect 40682 119200 40738 120000
rect 42246 119200 42302 120000
rect 43810 119200 43866 120000
rect 45374 119200 45430 120000
rect 46938 119200 46994 120000
rect 48502 119200 48558 120000
rect 50066 119200 50122 120000
rect 51630 119200 51686 120000
rect 53194 119200 53250 120000
rect 54758 119200 54814 120000
rect 56322 119200 56378 120000
rect 57886 119200 57942 120000
rect 59450 119200 59506 120000
rect 61014 119200 61070 120000
rect 62578 119200 62634 120000
rect 64142 119200 64198 120000
rect 65706 119200 65762 120000
rect 67270 119200 67326 120000
rect 68834 119200 68890 120000
rect 70398 119200 70454 120000
rect 71962 119200 72018 120000
rect 73526 119200 73582 120000
rect 75090 119200 75146 120000
rect 76654 119200 76710 120000
rect 78218 119200 78274 120000
rect 79782 119200 79838 120000
rect 81346 119200 81402 120000
rect 82910 119200 82966 120000
rect 84474 119200 84530 120000
rect 86038 119200 86094 120000
rect 87602 119200 87658 120000
rect 89166 119200 89222 120000
rect 90730 119200 90786 120000
rect 92294 119200 92350 120000
rect 93858 119200 93914 120000
rect 95422 119200 95478 120000
rect 96986 119200 97042 120000
rect 98550 119200 98606 120000
rect 100114 119200 100170 120000
rect 101678 119200 101734 120000
rect 103242 119200 103298 120000
rect 104806 119200 104862 120000
rect 106370 119200 106426 120000
rect 107934 119200 107990 120000
rect 109498 119200 109554 120000
rect 111062 119200 111118 120000
rect 112626 119200 112682 120000
rect 114190 119200 114246 120000
rect 115754 119200 115810 120000
rect 117318 119200 117374 120000
rect 118882 119200 118938 120000
rect 120446 119200 120502 120000
rect 122010 119200 122066 120000
rect 123574 119200 123630 120000
rect 125138 119200 125194 120000
rect 126702 119200 126758 120000
rect 128266 119200 128322 120000
rect 129830 119200 129886 120000
rect 131394 119200 131450 120000
rect 132958 119200 133014 120000
rect 134522 119200 134578 120000
rect 136086 119200 136142 120000
rect 137650 119200 137706 120000
rect 139214 119200 139270 120000
rect 140778 119200 140834 120000
rect 142342 119200 142398 120000
rect 143906 119200 143962 120000
rect 145470 119200 145526 120000
rect 147034 119200 147090 120000
rect 148598 119200 148654 120000
rect 150162 119200 150218 120000
rect 151726 119200 151782 120000
rect 153290 119200 153346 120000
rect 154854 119200 154910 120000
rect 156418 119200 156474 120000
rect 157982 119200 158038 120000
rect 159546 119200 159602 120000
rect 161110 119200 161166 120000
rect 162674 119200 162730 120000
rect 164238 119200 164294 120000
rect 165802 119200 165858 120000
rect 167366 119200 167422 120000
rect 168930 119200 168986 120000
rect 170494 119200 170550 120000
rect 172058 119200 172114 120000
rect 173622 119200 173678 120000
rect 175186 119200 175242 120000
rect 176750 119200 176806 120000
rect 178314 119200 178370 120000
rect 22006 0 22062 800
rect 22282 0 22338 800
rect 22558 0 22614 800
rect 22834 0 22890 800
rect 23110 0 23166 800
rect 23386 0 23442 800
rect 23662 0 23718 800
rect 23938 0 23994 800
rect 24214 0 24270 800
rect 24490 0 24546 800
rect 24766 0 24822 800
rect 25042 0 25098 800
rect 25318 0 25374 800
rect 25594 0 25650 800
rect 25870 0 25926 800
rect 26146 0 26202 800
rect 26422 0 26478 800
rect 26698 0 26754 800
rect 26974 0 27030 800
rect 27250 0 27306 800
rect 27526 0 27582 800
rect 27802 0 27858 800
rect 28078 0 28134 800
rect 28354 0 28410 800
rect 28630 0 28686 800
rect 28906 0 28962 800
rect 29182 0 29238 800
rect 29458 0 29514 800
rect 29734 0 29790 800
rect 30010 0 30066 800
rect 30286 0 30342 800
rect 30562 0 30618 800
rect 30838 0 30894 800
rect 31114 0 31170 800
rect 31390 0 31446 800
rect 31666 0 31722 800
rect 31942 0 31998 800
rect 32218 0 32274 800
rect 32494 0 32550 800
rect 32770 0 32826 800
rect 33046 0 33102 800
rect 33322 0 33378 800
rect 33598 0 33654 800
rect 33874 0 33930 800
rect 34150 0 34206 800
rect 34426 0 34482 800
rect 34702 0 34758 800
rect 34978 0 35034 800
rect 35254 0 35310 800
rect 35530 0 35586 800
rect 35806 0 35862 800
rect 36082 0 36138 800
rect 36358 0 36414 800
rect 36634 0 36690 800
rect 36910 0 36966 800
rect 37186 0 37242 800
rect 37462 0 37518 800
rect 37738 0 37794 800
rect 38014 0 38070 800
rect 38290 0 38346 800
rect 38566 0 38622 800
rect 38842 0 38898 800
rect 39118 0 39174 800
rect 39394 0 39450 800
rect 39670 0 39726 800
rect 39946 0 40002 800
rect 40222 0 40278 800
rect 40498 0 40554 800
rect 40774 0 40830 800
rect 41050 0 41106 800
rect 41326 0 41382 800
rect 41602 0 41658 800
rect 41878 0 41934 800
rect 42154 0 42210 800
rect 42430 0 42486 800
rect 42706 0 42762 800
rect 42982 0 43038 800
rect 43258 0 43314 800
rect 43534 0 43590 800
rect 43810 0 43866 800
rect 44086 0 44142 800
rect 44362 0 44418 800
rect 44638 0 44694 800
rect 44914 0 44970 800
rect 45190 0 45246 800
rect 45466 0 45522 800
rect 45742 0 45798 800
rect 46018 0 46074 800
rect 46294 0 46350 800
rect 46570 0 46626 800
rect 46846 0 46902 800
rect 47122 0 47178 800
rect 47398 0 47454 800
rect 47674 0 47730 800
rect 47950 0 48006 800
rect 48226 0 48282 800
rect 48502 0 48558 800
rect 48778 0 48834 800
rect 49054 0 49110 800
rect 49330 0 49386 800
rect 49606 0 49662 800
rect 49882 0 49938 800
rect 50158 0 50214 800
rect 50434 0 50490 800
rect 50710 0 50766 800
rect 50986 0 51042 800
rect 51262 0 51318 800
rect 51538 0 51594 800
rect 51814 0 51870 800
rect 52090 0 52146 800
rect 52366 0 52422 800
rect 52642 0 52698 800
rect 52918 0 52974 800
rect 53194 0 53250 800
rect 53470 0 53526 800
rect 53746 0 53802 800
rect 54022 0 54078 800
rect 54298 0 54354 800
rect 54574 0 54630 800
rect 54850 0 54906 800
rect 55126 0 55182 800
rect 55402 0 55458 800
rect 55678 0 55734 800
rect 55954 0 56010 800
rect 56230 0 56286 800
rect 56506 0 56562 800
rect 56782 0 56838 800
rect 57058 0 57114 800
rect 57334 0 57390 800
rect 57610 0 57666 800
rect 57886 0 57942 800
rect 58162 0 58218 800
rect 58438 0 58494 800
rect 58714 0 58770 800
rect 58990 0 59046 800
rect 59266 0 59322 800
rect 59542 0 59598 800
rect 59818 0 59874 800
rect 60094 0 60150 800
rect 60370 0 60426 800
rect 60646 0 60702 800
rect 60922 0 60978 800
rect 61198 0 61254 800
rect 61474 0 61530 800
rect 61750 0 61806 800
rect 62026 0 62082 800
rect 62302 0 62358 800
rect 62578 0 62634 800
rect 62854 0 62910 800
rect 63130 0 63186 800
rect 63406 0 63462 800
rect 63682 0 63738 800
rect 63958 0 64014 800
rect 64234 0 64290 800
rect 64510 0 64566 800
rect 64786 0 64842 800
rect 65062 0 65118 800
rect 65338 0 65394 800
rect 65614 0 65670 800
rect 65890 0 65946 800
rect 66166 0 66222 800
rect 66442 0 66498 800
rect 66718 0 66774 800
rect 66994 0 67050 800
rect 67270 0 67326 800
rect 67546 0 67602 800
rect 67822 0 67878 800
rect 68098 0 68154 800
rect 68374 0 68430 800
rect 68650 0 68706 800
rect 68926 0 68982 800
rect 69202 0 69258 800
rect 69478 0 69534 800
rect 69754 0 69810 800
rect 70030 0 70086 800
rect 70306 0 70362 800
rect 70582 0 70638 800
rect 70858 0 70914 800
rect 71134 0 71190 800
rect 71410 0 71466 800
rect 71686 0 71742 800
rect 71962 0 72018 800
rect 72238 0 72294 800
rect 72514 0 72570 800
rect 72790 0 72846 800
rect 73066 0 73122 800
rect 73342 0 73398 800
rect 73618 0 73674 800
rect 73894 0 73950 800
rect 74170 0 74226 800
rect 74446 0 74502 800
rect 74722 0 74778 800
rect 74998 0 75054 800
rect 75274 0 75330 800
rect 75550 0 75606 800
rect 75826 0 75882 800
rect 76102 0 76158 800
rect 76378 0 76434 800
rect 76654 0 76710 800
rect 76930 0 76986 800
rect 77206 0 77262 800
rect 77482 0 77538 800
rect 77758 0 77814 800
rect 78034 0 78090 800
rect 78310 0 78366 800
rect 78586 0 78642 800
rect 78862 0 78918 800
rect 79138 0 79194 800
rect 79414 0 79470 800
rect 79690 0 79746 800
rect 79966 0 80022 800
rect 80242 0 80298 800
rect 80518 0 80574 800
rect 80794 0 80850 800
rect 81070 0 81126 800
rect 81346 0 81402 800
rect 81622 0 81678 800
rect 81898 0 81954 800
rect 82174 0 82230 800
rect 82450 0 82506 800
rect 82726 0 82782 800
rect 83002 0 83058 800
rect 83278 0 83334 800
rect 83554 0 83610 800
rect 83830 0 83886 800
rect 84106 0 84162 800
rect 84382 0 84438 800
rect 84658 0 84714 800
rect 84934 0 84990 800
rect 85210 0 85266 800
rect 85486 0 85542 800
rect 85762 0 85818 800
rect 86038 0 86094 800
rect 86314 0 86370 800
rect 86590 0 86646 800
rect 86866 0 86922 800
rect 87142 0 87198 800
rect 87418 0 87474 800
rect 87694 0 87750 800
rect 87970 0 88026 800
rect 88246 0 88302 800
rect 88522 0 88578 800
rect 88798 0 88854 800
rect 89074 0 89130 800
rect 89350 0 89406 800
rect 89626 0 89682 800
rect 89902 0 89958 800
rect 90178 0 90234 800
rect 90454 0 90510 800
rect 90730 0 90786 800
rect 91006 0 91062 800
rect 91282 0 91338 800
rect 91558 0 91614 800
rect 91834 0 91890 800
rect 92110 0 92166 800
rect 92386 0 92442 800
rect 92662 0 92718 800
rect 92938 0 92994 800
rect 93214 0 93270 800
rect 93490 0 93546 800
rect 93766 0 93822 800
rect 94042 0 94098 800
rect 94318 0 94374 800
rect 94594 0 94650 800
rect 94870 0 94926 800
rect 95146 0 95202 800
rect 95422 0 95478 800
rect 95698 0 95754 800
rect 95974 0 96030 800
rect 96250 0 96306 800
rect 96526 0 96582 800
rect 96802 0 96858 800
rect 97078 0 97134 800
rect 97354 0 97410 800
rect 97630 0 97686 800
rect 97906 0 97962 800
rect 98182 0 98238 800
rect 98458 0 98514 800
rect 98734 0 98790 800
rect 99010 0 99066 800
rect 99286 0 99342 800
rect 99562 0 99618 800
rect 99838 0 99894 800
rect 100114 0 100170 800
rect 100390 0 100446 800
rect 100666 0 100722 800
rect 100942 0 100998 800
rect 101218 0 101274 800
rect 101494 0 101550 800
rect 101770 0 101826 800
rect 102046 0 102102 800
rect 102322 0 102378 800
rect 102598 0 102654 800
rect 102874 0 102930 800
rect 103150 0 103206 800
rect 103426 0 103482 800
rect 103702 0 103758 800
rect 103978 0 104034 800
rect 104254 0 104310 800
rect 104530 0 104586 800
rect 104806 0 104862 800
rect 105082 0 105138 800
rect 105358 0 105414 800
rect 105634 0 105690 800
rect 105910 0 105966 800
rect 106186 0 106242 800
rect 106462 0 106518 800
rect 106738 0 106794 800
rect 107014 0 107070 800
rect 107290 0 107346 800
rect 107566 0 107622 800
rect 107842 0 107898 800
rect 108118 0 108174 800
rect 108394 0 108450 800
rect 108670 0 108726 800
rect 108946 0 109002 800
rect 109222 0 109278 800
rect 109498 0 109554 800
rect 109774 0 109830 800
rect 110050 0 110106 800
rect 110326 0 110382 800
rect 110602 0 110658 800
rect 110878 0 110934 800
rect 111154 0 111210 800
rect 111430 0 111486 800
rect 111706 0 111762 800
rect 111982 0 112038 800
rect 112258 0 112314 800
rect 112534 0 112590 800
rect 112810 0 112866 800
rect 113086 0 113142 800
rect 113362 0 113418 800
rect 113638 0 113694 800
rect 113914 0 113970 800
rect 114190 0 114246 800
rect 114466 0 114522 800
rect 114742 0 114798 800
rect 115018 0 115074 800
rect 115294 0 115350 800
rect 115570 0 115626 800
rect 115846 0 115902 800
rect 116122 0 116178 800
rect 116398 0 116454 800
rect 116674 0 116730 800
rect 116950 0 117006 800
rect 117226 0 117282 800
rect 117502 0 117558 800
rect 117778 0 117834 800
rect 118054 0 118110 800
rect 118330 0 118386 800
rect 118606 0 118662 800
rect 118882 0 118938 800
rect 119158 0 119214 800
rect 119434 0 119490 800
rect 119710 0 119766 800
rect 119986 0 120042 800
rect 120262 0 120318 800
rect 120538 0 120594 800
rect 120814 0 120870 800
rect 121090 0 121146 800
rect 121366 0 121422 800
rect 121642 0 121698 800
rect 121918 0 121974 800
rect 122194 0 122250 800
rect 122470 0 122526 800
rect 122746 0 122802 800
rect 123022 0 123078 800
rect 123298 0 123354 800
rect 123574 0 123630 800
rect 123850 0 123906 800
rect 124126 0 124182 800
rect 124402 0 124458 800
rect 124678 0 124734 800
rect 124954 0 125010 800
rect 125230 0 125286 800
rect 125506 0 125562 800
rect 125782 0 125838 800
rect 126058 0 126114 800
rect 126334 0 126390 800
rect 126610 0 126666 800
rect 126886 0 126942 800
rect 127162 0 127218 800
rect 127438 0 127494 800
rect 127714 0 127770 800
rect 127990 0 128046 800
rect 128266 0 128322 800
rect 128542 0 128598 800
rect 128818 0 128874 800
rect 129094 0 129150 800
rect 129370 0 129426 800
rect 129646 0 129702 800
rect 129922 0 129978 800
rect 130198 0 130254 800
rect 130474 0 130530 800
rect 130750 0 130806 800
rect 131026 0 131082 800
rect 131302 0 131358 800
rect 131578 0 131634 800
rect 131854 0 131910 800
rect 132130 0 132186 800
rect 132406 0 132462 800
rect 132682 0 132738 800
rect 132958 0 133014 800
rect 133234 0 133290 800
rect 133510 0 133566 800
rect 133786 0 133842 800
rect 134062 0 134118 800
rect 134338 0 134394 800
rect 134614 0 134670 800
rect 134890 0 134946 800
rect 135166 0 135222 800
rect 135442 0 135498 800
rect 135718 0 135774 800
rect 135994 0 136050 800
rect 136270 0 136326 800
rect 136546 0 136602 800
rect 136822 0 136878 800
rect 137098 0 137154 800
rect 137374 0 137430 800
rect 137650 0 137706 800
rect 137926 0 137982 800
rect 138202 0 138258 800
rect 138478 0 138534 800
rect 138754 0 138810 800
rect 139030 0 139086 800
rect 139306 0 139362 800
rect 139582 0 139638 800
rect 139858 0 139914 800
rect 140134 0 140190 800
rect 140410 0 140466 800
rect 140686 0 140742 800
rect 140962 0 141018 800
rect 141238 0 141294 800
rect 141514 0 141570 800
rect 141790 0 141846 800
rect 142066 0 142122 800
rect 142342 0 142398 800
rect 142618 0 142674 800
rect 142894 0 142950 800
rect 143170 0 143226 800
rect 143446 0 143502 800
rect 143722 0 143778 800
rect 143998 0 144054 800
rect 144274 0 144330 800
rect 144550 0 144606 800
rect 144826 0 144882 800
rect 145102 0 145158 800
rect 145378 0 145434 800
rect 145654 0 145710 800
rect 145930 0 145986 800
rect 146206 0 146262 800
rect 146482 0 146538 800
rect 146758 0 146814 800
rect 147034 0 147090 800
rect 147310 0 147366 800
rect 147586 0 147642 800
rect 147862 0 147918 800
rect 148138 0 148194 800
rect 148414 0 148470 800
rect 148690 0 148746 800
rect 148966 0 149022 800
rect 149242 0 149298 800
rect 149518 0 149574 800
rect 149794 0 149850 800
rect 150070 0 150126 800
rect 150346 0 150402 800
rect 150622 0 150678 800
rect 150898 0 150954 800
rect 151174 0 151230 800
rect 151450 0 151506 800
rect 151726 0 151782 800
rect 152002 0 152058 800
rect 152278 0 152334 800
rect 152554 0 152610 800
rect 152830 0 152886 800
rect 153106 0 153162 800
rect 153382 0 153438 800
rect 153658 0 153714 800
rect 153934 0 153990 800
rect 154210 0 154266 800
rect 154486 0 154542 800
rect 154762 0 154818 800
rect 155038 0 155094 800
rect 155314 0 155370 800
rect 155590 0 155646 800
rect 155866 0 155922 800
rect 156142 0 156198 800
rect 156418 0 156474 800
rect 156694 0 156750 800
rect 156970 0 157026 800
rect 157246 0 157302 800
rect 157522 0 157578 800
rect 157798 0 157854 800
<< obsm2 >>
rect 3258 119144 4654 119354
rect 4822 119144 6218 119354
rect 6386 119144 7782 119354
rect 7950 119144 9346 119354
rect 9514 119144 10910 119354
rect 11078 119144 12474 119354
rect 12642 119144 14038 119354
rect 14206 119144 15602 119354
rect 15770 119144 17166 119354
rect 17334 119144 18730 119354
rect 18898 119144 20294 119354
rect 20462 119144 21858 119354
rect 22026 119144 23422 119354
rect 23590 119144 24986 119354
rect 25154 119144 26550 119354
rect 26718 119144 28114 119354
rect 28282 119144 29678 119354
rect 29846 119144 31242 119354
rect 31410 119144 32806 119354
rect 32974 119144 34370 119354
rect 34538 119144 35934 119354
rect 36102 119144 37498 119354
rect 37666 119144 39062 119354
rect 39230 119144 40626 119354
rect 40794 119144 42190 119354
rect 42358 119144 43754 119354
rect 43922 119144 45318 119354
rect 45486 119144 46882 119354
rect 47050 119144 48446 119354
rect 48614 119144 50010 119354
rect 50178 119144 51574 119354
rect 51742 119144 53138 119354
rect 53306 119144 54702 119354
rect 54870 119144 56266 119354
rect 56434 119144 57830 119354
rect 57998 119144 59394 119354
rect 59562 119144 60958 119354
rect 61126 119144 62522 119354
rect 62690 119144 64086 119354
rect 64254 119144 65650 119354
rect 65818 119144 67214 119354
rect 67382 119144 68778 119354
rect 68946 119144 70342 119354
rect 70510 119144 71906 119354
rect 72074 119144 73470 119354
rect 73638 119144 75034 119354
rect 75202 119144 76598 119354
rect 76766 119144 78162 119354
rect 78330 119144 79726 119354
rect 79894 119144 81290 119354
rect 81458 119144 82854 119354
rect 83022 119144 84418 119354
rect 84586 119144 85982 119354
rect 86150 119144 87546 119354
rect 87714 119144 89110 119354
rect 89278 119144 90674 119354
rect 90842 119144 92238 119354
rect 92406 119144 93802 119354
rect 93970 119144 95366 119354
rect 95534 119144 96930 119354
rect 97098 119144 98494 119354
rect 98662 119144 100058 119354
rect 100226 119144 101622 119354
rect 101790 119144 103186 119354
rect 103354 119144 104750 119354
rect 104918 119144 106314 119354
rect 106482 119144 107878 119354
rect 108046 119144 109442 119354
rect 109610 119144 111006 119354
rect 111174 119144 112570 119354
rect 112738 119144 114134 119354
rect 114302 119144 115698 119354
rect 115866 119144 117262 119354
rect 117430 119144 118826 119354
rect 118994 119144 120390 119354
rect 120558 119144 121954 119354
rect 122122 119144 123518 119354
rect 123686 119144 125082 119354
rect 125250 119144 126646 119354
rect 126814 119144 128210 119354
rect 128378 119144 129774 119354
rect 129942 119144 131338 119354
rect 131506 119144 132902 119354
rect 133070 119144 134466 119354
rect 134634 119144 136030 119354
rect 136198 119144 137594 119354
rect 137762 119144 139158 119354
rect 139326 119144 140722 119354
rect 140890 119144 142286 119354
rect 142454 119144 143850 119354
rect 144018 119144 145414 119354
rect 145582 119144 146978 119354
rect 147146 119144 148542 119354
rect 148710 119144 150106 119354
rect 150274 119144 151670 119354
rect 151838 119144 153234 119354
rect 153402 119144 154798 119354
rect 154966 119144 156362 119354
rect 156530 119144 157926 119354
rect 158094 119144 159490 119354
rect 159658 119144 161054 119354
rect 161222 119144 162618 119354
rect 162786 119144 164182 119354
rect 164350 119144 165746 119354
rect 165914 119144 167310 119354
rect 167478 119144 168874 119354
rect 169042 119144 170438 119354
rect 170606 119144 172002 119354
rect 172170 119144 173566 119354
rect 173734 119144 175130 119354
rect 175298 119144 176694 119354
rect 176862 119144 178258 119354
rect 3202 856 178368 119144
rect 3202 800 21950 856
rect 22118 800 22226 856
rect 22394 800 22502 856
rect 22670 800 22778 856
rect 22946 800 23054 856
rect 23222 800 23330 856
rect 23498 800 23606 856
rect 23774 800 23882 856
rect 24050 800 24158 856
rect 24326 800 24434 856
rect 24602 800 24710 856
rect 24878 800 24986 856
rect 25154 800 25262 856
rect 25430 800 25538 856
rect 25706 800 25814 856
rect 25982 800 26090 856
rect 26258 800 26366 856
rect 26534 800 26642 856
rect 26810 800 26918 856
rect 27086 800 27194 856
rect 27362 800 27470 856
rect 27638 800 27746 856
rect 27914 800 28022 856
rect 28190 800 28298 856
rect 28466 800 28574 856
rect 28742 800 28850 856
rect 29018 800 29126 856
rect 29294 800 29402 856
rect 29570 800 29678 856
rect 29846 800 29954 856
rect 30122 800 30230 856
rect 30398 800 30506 856
rect 30674 800 30782 856
rect 30950 800 31058 856
rect 31226 800 31334 856
rect 31502 800 31610 856
rect 31778 800 31886 856
rect 32054 800 32162 856
rect 32330 800 32438 856
rect 32606 800 32714 856
rect 32882 800 32990 856
rect 33158 800 33266 856
rect 33434 800 33542 856
rect 33710 800 33818 856
rect 33986 800 34094 856
rect 34262 800 34370 856
rect 34538 800 34646 856
rect 34814 800 34922 856
rect 35090 800 35198 856
rect 35366 800 35474 856
rect 35642 800 35750 856
rect 35918 800 36026 856
rect 36194 800 36302 856
rect 36470 800 36578 856
rect 36746 800 36854 856
rect 37022 800 37130 856
rect 37298 800 37406 856
rect 37574 800 37682 856
rect 37850 800 37958 856
rect 38126 800 38234 856
rect 38402 800 38510 856
rect 38678 800 38786 856
rect 38954 800 39062 856
rect 39230 800 39338 856
rect 39506 800 39614 856
rect 39782 800 39890 856
rect 40058 800 40166 856
rect 40334 800 40442 856
rect 40610 800 40718 856
rect 40886 800 40994 856
rect 41162 800 41270 856
rect 41438 800 41546 856
rect 41714 800 41822 856
rect 41990 800 42098 856
rect 42266 800 42374 856
rect 42542 800 42650 856
rect 42818 800 42926 856
rect 43094 800 43202 856
rect 43370 800 43478 856
rect 43646 800 43754 856
rect 43922 800 44030 856
rect 44198 800 44306 856
rect 44474 800 44582 856
rect 44750 800 44858 856
rect 45026 800 45134 856
rect 45302 800 45410 856
rect 45578 800 45686 856
rect 45854 800 45962 856
rect 46130 800 46238 856
rect 46406 800 46514 856
rect 46682 800 46790 856
rect 46958 800 47066 856
rect 47234 800 47342 856
rect 47510 800 47618 856
rect 47786 800 47894 856
rect 48062 800 48170 856
rect 48338 800 48446 856
rect 48614 800 48722 856
rect 48890 800 48998 856
rect 49166 800 49274 856
rect 49442 800 49550 856
rect 49718 800 49826 856
rect 49994 800 50102 856
rect 50270 800 50378 856
rect 50546 800 50654 856
rect 50822 800 50930 856
rect 51098 800 51206 856
rect 51374 800 51482 856
rect 51650 800 51758 856
rect 51926 800 52034 856
rect 52202 800 52310 856
rect 52478 800 52586 856
rect 52754 800 52862 856
rect 53030 800 53138 856
rect 53306 800 53414 856
rect 53582 800 53690 856
rect 53858 800 53966 856
rect 54134 800 54242 856
rect 54410 800 54518 856
rect 54686 800 54794 856
rect 54962 800 55070 856
rect 55238 800 55346 856
rect 55514 800 55622 856
rect 55790 800 55898 856
rect 56066 800 56174 856
rect 56342 800 56450 856
rect 56618 800 56726 856
rect 56894 800 57002 856
rect 57170 800 57278 856
rect 57446 800 57554 856
rect 57722 800 57830 856
rect 57998 800 58106 856
rect 58274 800 58382 856
rect 58550 800 58658 856
rect 58826 800 58934 856
rect 59102 800 59210 856
rect 59378 800 59486 856
rect 59654 800 59762 856
rect 59930 800 60038 856
rect 60206 800 60314 856
rect 60482 800 60590 856
rect 60758 800 60866 856
rect 61034 800 61142 856
rect 61310 800 61418 856
rect 61586 800 61694 856
rect 61862 800 61970 856
rect 62138 800 62246 856
rect 62414 800 62522 856
rect 62690 800 62798 856
rect 62966 800 63074 856
rect 63242 800 63350 856
rect 63518 800 63626 856
rect 63794 800 63902 856
rect 64070 800 64178 856
rect 64346 800 64454 856
rect 64622 800 64730 856
rect 64898 800 65006 856
rect 65174 800 65282 856
rect 65450 800 65558 856
rect 65726 800 65834 856
rect 66002 800 66110 856
rect 66278 800 66386 856
rect 66554 800 66662 856
rect 66830 800 66938 856
rect 67106 800 67214 856
rect 67382 800 67490 856
rect 67658 800 67766 856
rect 67934 800 68042 856
rect 68210 800 68318 856
rect 68486 800 68594 856
rect 68762 800 68870 856
rect 69038 800 69146 856
rect 69314 800 69422 856
rect 69590 800 69698 856
rect 69866 800 69974 856
rect 70142 800 70250 856
rect 70418 800 70526 856
rect 70694 800 70802 856
rect 70970 800 71078 856
rect 71246 800 71354 856
rect 71522 800 71630 856
rect 71798 800 71906 856
rect 72074 800 72182 856
rect 72350 800 72458 856
rect 72626 800 72734 856
rect 72902 800 73010 856
rect 73178 800 73286 856
rect 73454 800 73562 856
rect 73730 800 73838 856
rect 74006 800 74114 856
rect 74282 800 74390 856
rect 74558 800 74666 856
rect 74834 800 74942 856
rect 75110 800 75218 856
rect 75386 800 75494 856
rect 75662 800 75770 856
rect 75938 800 76046 856
rect 76214 800 76322 856
rect 76490 800 76598 856
rect 76766 800 76874 856
rect 77042 800 77150 856
rect 77318 800 77426 856
rect 77594 800 77702 856
rect 77870 800 77978 856
rect 78146 800 78254 856
rect 78422 800 78530 856
rect 78698 800 78806 856
rect 78974 800 79082 856
rect 79250 800 79358 856
rect 79526 800 79634 856
rect 79802 800 79910 856
rect 80078 800 80186 856
rect 80354 800 80462 856
rect 80630 800 80738 856
rect 80906 800 81014 856
rect 81182 800 81290 856
rect 81458 800 81566 856
rect 81734 800 81842 856
rect 82010 800 82118 856
rect 82286 800 82394 856
rect 82562 800 82670 856
rect 82838 800 82946 856
rect 83114 800 83222 856
rect 83390 800 83498 856
rect 83666 800 83774 856
rect 83942 800 84050 856
rect 84218 800 84326 856
rect 84494 800 84602 856
rect 84770 800 84878 856
rect 85046 800 85154 856
rect 85322 800 85430 856
rect 85598 800 85706 856
rect 85874 800 85982 856
rect 86150 800 86258 856
rect 86426 800 86534 856
rect 86702 800 86810 856
rect 86978 800 87086 856
rect 87254 800 87362 856
rect 87530 800 87638 856
rect 87806 800 87914 856
rect 88082 800 88190 856
rect 88358 800 88466 856
rect 88634 800 88742 856
rect 88910 800 89018 856
rect 89186 800 89294 856
rect 89462 800 89570 856
rect 89738 800 89846 856
rect 90014 800 90122 856
rect 90290 800 90398 856
rect 90566 800 90674 856
rect 90842 800 90950 856
rect 91118 800 91226 856
rect 91394 800 91502 856
rect 91670 800 91778 856
rect 91946 800 92054 856
rect 92222 800 92330 856
rect 92498 800 92606 856
rect 92774 800 92882 856
rect 93050 800 93158 856
rect 93326 800 93434 856
rect 93602 800 93710 856
rect 93878 800 93986 856
rect 94154 800 94262 856
rect 94430 800 94538 856
rect 94706 800 94814 856
rect 94982 800 95090 856
rect 95258 800 95366 856
rect 95534 800 95642 856
rect 95810 800 95918 856
rect 96086 800 96194 856
rect 96362 800 96470 856
rect 96638 800 96746 856
rect 96914 800 97022 856
rect 97190 800 97298 856
rect 97466 800 97574 856
rect 97742 800 97850 856
rect 98018 800 98126 856
rect 98294 800 98402 856
rect 98570 800 98678 856
rect 98846 800 98954 856
rect 99122 800 99230 856
rect 99398 800 99506 856
rect 99674 800 99782 856
rect 99950 800 100058 856
rect 100226 800 100334 856
rect 100502 800 100610 856
rect 100778 800 100886 856
rect 101054 800 101162 856
rect 101330 800 101438 856
rect 101606 800 101714 856
rect 101882 800 101990 856
rect 102158 800 102266 856
rect 102434 800 102542 856
rect 102710 800 102818 856
rect 102986 800 103094 856
rect 103262 800 103370 856
rect 103538 800 103646 856
rect 103814 800 103922 856
rect 104090 800 104198 856
rect 104366 800 104474 856
rect 104642 800 104750 856
rect 104918 800 105026 856
rect 105194 800 105302 856
rect 105470 800 105578 856
rect 105746 800 105854 856
rect 106022 800 106130 856
rect 106298 800 106406 856
rect 106574 800 106682 856
rect 106850 800 106958 856
rect 107126 800 107234 856
rect 107402 800 107510 856
rect 107678 800 107786 856
rect 107954 800 108062 856
rect 108230 800 108338 856
rect 108506 800 108614 856
rect 108782 800 108890 856
rect 109058 800 109166 856
rect 109334 800 109442 856
rect 109610 800 109718 856
rect 109886 800 109994 856
rect 110162 800 110270 856
rect 110438 800 110546 856
rect 110714 800 110822 856
rect 110990 800 111098 856
rect 111266 800 111374 856
rect 111542 800 111650 856
rect 111818 800 111926 856
rect 112094 800 112202 856
rect 112370 800 112478 856
rect 112646 800 112754 856
rect 112922 800 113030 856
rect 113198 800 113306 856
rect 113474 800 113582 856
rect 113750 800 113858 856
rect 114026 800 114134 856
rect 114302 800 114410 856
rect 114578 800 114686 856
rect 114854 800 114962 856
rect 115130 800 115238 856
rect 115406 800 115514 856
rect 115682 800 115790 856
rect 115958 800 116066 856
rect 116234 800 116342 856
rect 116510 800 116618 856
rect 116786 800 116894 856
rect 117062 800 117170 856
rect 117338 800 117446 856
rect 117614 800 117722 856
rect 117890 800 117998 856
rect 118166 800 118274 856
rect 118442 800 118550 856
rect 118718 800 118826 856
rect 118994 800 119102 856
rect 119270 800 119378 856
rect 119546 800 119654 856
rect 119822 800 119930 856
rect 120098 800 120206 856
rect 120374 800 120482 856
rect 120650 800 120758 856
rect 120926 800 121034 856
rect 121202 800 121310 856
rect 121478 800 121586 856
rect 121754 800 121862 856
rect 122030 800 122138 856
rect 122306 800 122414 856
rect 122582 800 122690 856
rect 122858 800 122966 856
rect 123134 800 123242 856
rect 123410 800 123518 856
rect 123686 800 123794 856
rect 123962 800 124070 856
rect 124238 800 124346 856
rect 124514 800 124622 856
rect 124790 800 124898 856
rect 125066 800 125174 856
rect 125342 800 125450 856
rect 125618 800 125726 856
rect 125894 800 126002 856
rect 126170 800 126278 856
rect 126446 800 126554 856
rect 126722 800 126830 856
rect 126998 800 127106 856
rect 127274 800 127382 856
rect 127550 800 127658 856
rect 127826 800 127934 856
rect 128102 800 128210 856
rect 128378 800 128486 856
rect 128654 800 128762 856
rect 128930 800 129038 856
rect 129206 800 129314 856
rect 129482 800 129590 856
rect 129758 800 129866 856
rect 130034 800 130142 856
rect 130310 800 130418 856
rect 130586 800 130694 856
rect 130862 800 130970 856
rect 131138 800 131246 856
rect 131414 800 131522 856
rect 131690 800 131798 856
rect 131966 800 132074 856
rect 132242 800 132350 856
rect 132518 800 132626 856
rect 132794 800 132902 856
rect 133070 800 133178 856
rect 133346 800 133454 856
rect 133622 800 133730 856
rect 133898 800 134006 856
rect 134174 800 134282 856
rect 134450 800 134558 856
rect 134726 800 134834 856
rect 135002 800 135110 856
rect 135278 800 135386 856
rect 135554 800 135662 856
rect 135830 800 135938 856
rect 136106 800 136214 856
rect 136382 800 136490 856
rect 136658 800 136766 856
rect 136934 800 137042 856
rect 137210 800 137318 856
rect 137486 800 137594 856
rect 137762 800 137870 856
rect 138038 800 138146 856
rect 138314 800 138422 856
rect 138590 800 138698 856
rect 138866 800 138974 856
rect 139142 800 139250 856
rect 139418 800 139526 856
rect 139694 800 139802 856
rect 139970 800 140078 856
rect 140246 800 140354 856
rect 140522 800 140630 856
rect 140798 800 140906 856
rect 141074 800 141182 856
rect 141350 800 141458 856
rect 141626 800 141734 856
rect 141902 800 142010 856
rect 142178 800 142286 856
rect 142454 800 142562 856
rect 142730 800 142838 856
rect 143006 800 143114 856
rect 143282 800 143390 856
rect 143558 800 143666 856
rect 143834 800 143942 856
rect 144110 800 144218 856
rect 144386 800 144494 856
rect 144662 800 144770 856
rect 144938 800 145046 856
rect 145214 800 145322 856
rect 145490 800 145598 856
rect 145766 800 145874 856
rect 146042 800 146150 856
rect 146318 800 146426 856
rect 146594 800 146702 856
rect 146870 800 146978 856
rect 147146 800 147254 856
rect 147422 800 147530 856
rect 147698 800 147806 856
rect 147974 800 148082 856
rect 148250 800 148358 856
rect 148526 800 148634 856
rect 148802 800 148910 856
rect 149078 800 149186 856
rect 149354 800 149462 856
rect 149630 800 149738 856
rect 149906 800 150014 856
rect 150182 800 150290 856
rect 150458 800 150566 856
rect 150734 800 150842 856
rect 151010 800 151118 856
rect 151286 800 151394 856
rect 151562 800 151670 856
rect 151838 800 151946 856
rect 152114 800 152222 856
rect 152390 800 152498 856
rect 152666 800 152774 856
rect 152942 800 153050 856
rect 153218 800 153326 856
rect 153494 800 153602 856
rect 153770 800 153878 856
rect 154046 800 154154 856
rect 154322 800 154430 856
rect 154598 800 154706 856
rect 154874 800 154982 856
rect 155150 800 155258 856
rect 155426 800 155534 856
rect 155702 800 155810 856
rect 155978 800 156086 856
rect 156254 800 156362 856
rect 156530 800 156638 856
rect 156806 800 156914 856
rect 157082 800 157190 856
rect 157358 800 157466 856
rect 157634 800 157742 856
rect 157910 800 178368 856
<< obsm3 >>
rect 4210 2143 173486 117537
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< labels >>
rlabel metal2 s 1582 119200 1638 120000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 48502 119200 48558 120000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 53194 119200 53250 120000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 57886 119200 57942 120000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 62578 119200 62634 120000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 67270 119200 67326 120000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 71962 119200 72018 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 76654 119200 76710 120000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 81346 119200 81402 120000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 86038 119200 86094 120000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 90730 119200 90786 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 6274 119200 6330 120000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 95422 119200 95478 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 100114 119200 100170 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 104806 119200 104862 120000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 109498 119200 109554 120000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 114190 119200 114246 120000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 118882 119200 118938 120000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 123574 119200 123630 120000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 128266 119200 128322 120000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 132958 119200 133014 120000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 137650 119200 137706 120000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 10966 119200 11022 120000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 142342 119200 142398 120000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 147034 119200 147090 120000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 151726 119200 151782 120000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 156418 119200 156474 120000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 161110 119200 161166 120000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 165802 119200 165858 120000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 170494 119200 170550 120000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 175186 119200 175242 120000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 15658 119200 15714 120000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 20350 119200 20406 120000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 25042 119200 25098 120000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 29734 119200 29790 120000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 34426 119200 34482 120000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 39118 119200 39174 120000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 43810 119200 43866 120000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3146 119200 3202 120000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 50066 119200 50122 120000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 54758 119200 54814 120000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 59450 119200 59506 120000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 64142 119200 64198 120000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 68834 119200 68890 120000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 73526 119200 73582 120000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 78218 119200 78274 120000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 82910 119200 82966 120000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 87602 119200 87658 120000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 92294 119200 92350 120000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7838 119200 7894 120000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 96986 119200 97042 120000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 101678 119200 101734 120000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 106370 119200 106426 120000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 111062 119200 111118 120000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 115754 119200 115810 120000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 120446 119200 120502 120000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 125138 119200 125194 120000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 129830 119200 129886 120000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 134522 119200 134578 120000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 139214 119200 139270 120000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 12530 119200 12586 120000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 143906 119200 143962 120000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 148598 119200 148654 120000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 153290 119200 153346 120000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 157982 119200 158038 120000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 162674 119200 162730 120000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 167366 119200 167422 120000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 172058 119200 172114 120000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 176750 119200 176806 120000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 17222 119200 17278 120000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 21914 119200 21970 120000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 26606 119200 26662 120000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 31298 119200 31354 120000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 35990 119200 36046 120000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 40682 119200 40738 120000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 45374 119200 45430 120000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4710 119200 4766 120000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 51630 119200 51686 120000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 56322 119200 56378 120000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 61014 119200 61070 120000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 65706 119200 65762 120000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 70398 119200 70454 120000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 75090 119200 75146 120000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 79782 119200 79838 120000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 84474 119200 84530 120000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 89166 119200 89222 120000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 93858 119200 93914 120000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 9402 119200 9458 120000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 98550 119200 98606 120000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 103242 119200 103298 120000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 107934 119200 107990 120000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 112626 119200 112682 120000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 117318 119200 117374 120000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 122010 119200 122066 120000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 126702 119200 126758 120000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 131394 119200 131450 120000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 136086 119200 136142 120000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 140778 119200 140834 120000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 14094 119200 14150 120000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 145470 119200 145526 120000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 150162 119200 150218 120000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 154854 119200 154910 120000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 159546 119200 159602 120000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 164238 119200 164294 120000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 168930 119200 168986 120000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 173622 119200 173678 120000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 178314 119200 178370 120000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 18786 119200 18842 120000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 23478 119200 23534 120000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 28170 119200 28226 120000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 32862 119200 32918 120000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 37554 119200 37610 120000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 42246 119200 42302 120000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 46938 119200 46994 120000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 157246 0 157302 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 157522 0 157578 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 157798 0 157854 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 135718 0 135774 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 139030 0 139086 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 139858 0 139914 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 140686 0 140742 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 143998 0 144054 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 145654 0 145710 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 146482 0 146538 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 147310 0 147366 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 148966 0 149022 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 149794 0 149850 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 151450 0 151506 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 152278 0 152334 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 153106 0 153162 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 154762 0 154818 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 156418 0 156474 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 91834 0 91890 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 108394 0 108450 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 118330 0 118386 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 119986 0 120042 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 122470 0 122526 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 123298 0 123354 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 127438 0 127494 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 128266 0 128322 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 132406 0 132462 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 133234 0 133290 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 134338 0 134394 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 135166 0 135222 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 135994 0 136050 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 136822 0 136878 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 137650 0 137706 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 138478 0 138534 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 139306 0 139362 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 140134 0 140190 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 140962 0 141018 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 141790 0 141846 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 142618 0 142674 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 143446 0 143502 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 144274 0 144330 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 145102 0 145158 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 145930 0 145986 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 146758 0 146814 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 147586 0 147642 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 148414 0 148470 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 149242 0 149298 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 150070 0 150126 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 150898 0 150954 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 151726 0 151782 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 152554 0 152610 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 153382 0 153438 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 154210 0 154266 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 155038 0 155094 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 156694 0 156750 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 61474 0 61530 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 67270 0 67326 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 52366 0 52422 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 68098 0 68154 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 70582 0 70638 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 71410 0 71466 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 72238 0 72294 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 73066 0 73122 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 73894 0 73950 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 53194 0 53250 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 77206 0 77262 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 78034 0 78090 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 78862 0 78918 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 79690 0 79746 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 81346 0 81402 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 82174 0 82230 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 83002 0 83058 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 83830 0 83886 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 85486 0 85542 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 87142 0 87198 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 87970 0 88026 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 89626 0 89682 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 90454 0 90510 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 91282 0 91338 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 54850 0 54906 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 92938 0 92994 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 93766 0 93822 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 94594 0 94650 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 95422 0 95478 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 97078 0 97134 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 98734 0 98790 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 99562 0 99618 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 100390 0 100446 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 55678 0 55734 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 101218 0 101274 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 102046 0 102102 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 102874 0 102930 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 103702 0 103758 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 104530 0 104586 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 105358 0 105414 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 106186 0 106242 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 107014 0 107070 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 107842 0 107898 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 108670 0 108726 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 56506 0 56562 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 110326 0 110382 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 111154 0 111210 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 112810 0 112866 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 114466 0 114522 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 115294 0 115350 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 116122 0 116178 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 116950 0 117006 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 117778 0 117834 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 118606 0 118662 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 119434 0 119490 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 120262 0 120318 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 122746 0 122802 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 123574 0 123630 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 124402 0 124458 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 125230 0 125286 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 126058 0 126114 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 126886 0 126942 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 127714 0 127770 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 128542 0 128598 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 129370 0 129426 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 130198 0 130254 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 131026 0 131082 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 131854 0 131910 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 132682 0 132738 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 133510 0 133566 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 135442 0 135498 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 139582 0 139638 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 142066 0 142122 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 142894 0 142950 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 144550 0 144606 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 145378 0 145434 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 147862 0 147918 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 150346 0 150402 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 152830 0 152886 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 154486 0 154542 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 155314 0 155370 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 156142 0 156198 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 122194 0 122250 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 132130 0 132186 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 22006 0 22062 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 37738 0 37794 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 39394 0 39450 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5789836
string GDS_FILE /home/ProgramFiles/16-bit-Brent-Kung-Adder-IC-Design/openlane/user_proj_example/runs/22_11_14_15_24/results/signoff/user_proj_example.magic.gds
string GDS_START 58840
<< end >>

